/////////////////////////////////////////////////////////////
//                                                         //
//              School of Software of SJTU                 //
//                                                         //
/////////////////////////////////////////////////////////////

module sc_computer(resetn, clock, mem_clk, pc, inst, aluout, memout, imem_clk, dmem_clk);
	input         resetn, clock, mem_clk;
	output [31:0] pc, inst, aluout, memout;
	output        imem_clk, dmem_clk;
	wire   [31:0] data;
	wire          wmem;

	sc_cpu cpu(clock, resetn, inst, memout, pc, wmem, aluout, data); // CPU module.
	sc_instmem imem(pc, inst, clock, mem_clk, imem_clk); // Instruction memory.
	sc_datamem dmem(aluout, data, memout, wmem, clock, mem_clk, dmem_clk); // Data memory.
endmodule
